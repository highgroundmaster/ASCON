`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/26/2023 05:58:13 PM
// Design Name: 
// Module Name: linear
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module linear(
    input [319:0] x,
    output [319:0] y
    );
    
  assign y[63:0] = x[63:0] ^ {x[(7-1):0], x[63:7]} ^ {x[(41-1):0], x[63:41]};
  assign y[127:64] = x[127:64] ^ {x[(64 + 10 - 1) :64], x[127: (64 + 10)]} ^ {x[(64 + 17 - 1):64], x[127:(64 + 17)]};
  assign y[191:128] = x[191:128] ^ {x[128], x[191:129]} ^ {x[(128 + 6 - 1):128], x[191:(128 + 6)]};
  assign y[255:192] = x[255:192] ^ {x[(192 + 61 -1):192], x[255:(192 + 61)]} ^ {x[(192 + 39 -1):192], x[255:(192 + 39)]};
  assign y[319:256] = x[319:256] ^ {x[(256 + 19 -1):256], x[319:(256+19)]} ^ {x[(256 + 28 -1):256], x[319:(256+28)]};

endmodule
